package env_pkg;

   `include "uvm_macros.svh"
   import uvm_pkg::*;

   
   `include "monitor.svh"
   `include "driver.svh"
   `include "sequencer.svh"

   `include "agent.svh"
   `include "env.svh"

endpackage

