package test_pkg;

   `include "uvm_macros.svh"
   import uvm_pkg::*;

   
   `include "base_test.svh"
   `include "sample_test.svh"

endpackage

